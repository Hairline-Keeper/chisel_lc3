`define RAMWIDTH 16

module RAMHelper(
    input                   clka,
    input                   ena,
    input                   wea,
    input   [`RAMWIDTH-1:0] addra,
    input   [`RAMWIDTH-1:0] dina,
    output  [`RAMWIDTH-1:0] douta

);

endmodule